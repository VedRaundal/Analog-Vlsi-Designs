module Alphabet_Gen(
    input  [5:0] D,
    input  [2:0] S,
    output reg [4:0] Alphabet
);

always @(*) begin
    case ({D, S})
        {6'd1, 3'd0}, {6'd1, 3'd1}, {6'd1, 3'd2}, {6'd1, 3'd3}, {6'd1, 3'd4}, {6'd1, 3'd5}:
            Alphabet = 5'd1;
        {6'd2, 3'd0}, {6'd2, 3'd1}, {6'd2, 3'd2}, {6'd2, 3'd3}, {6'd2, 3'd4}, {6'd2, 3'd5}:
            Alphabet = 5'd2;
        {6'd3, 3'd0}, {6'd3, 3'd1}, {6'd3, 3'd2}, {6'd3, 3'd3}, {6'd3, 3'd4}, {6'd3, 3'd5}:
            Alphabet = 5'd3;
        {6'd4, 3'd0}, {6'd4, 3'd1}, {6'd4, 3'd2}, {6'd4, 3'd3}, {6'd4, 3'd4}, {6'd4, 3'd5}:
            Alphabet = 5'd4;
        {6'd5, 3'd0}, {6'd5, 3'd1}, {6'd5, 3'd2}, {6'd5, 3'd3}, {6'd5, 3'd4}, {6'd5, 3'd5}:
            Alphabet = 5'd5;

        {6'd6, 3'd0}, {6'd6, 3'd1}, {6'd6, 3'd2}, {6'd6, 3'd3}, {6'd6, 3'd4}, {6'd6, 3'd5}:
            Alphabet = 5'd6;

        {6'd7, 3'd0},{6'd7, 3'd1}, {6'd7, 3'd2}, {6'd7, 3'd3}, {6'd7, 3'd4}, {6'd7, 3'd5}:
            Alphabet = 5'd6;
           

        {6'd8, 3'd0}, {6'd9, 3'd0}, {6'd10, 3'd0}:
            Alphabet = 5'd7;
        {6'd8, 3'd1}, {6'd8, 3'd2}, {6'd8, 3'd3}, {6'd8, 3'd4}, {6'd8, 3'd5},
        {6'd9, 3'd1}, {6'd9, 3'd2}, {6'd9, 3'd3}, {6'd9, 3'd4}, {6'd9, 3'd5},
        {6'd10, 3'd1}, {6'd10, 3'd2}, {6'd10, 3'd3}, {6'd10, 3'd4}, {6'd10, 3'd5}:
            Alphabet = 5'd8;

        {6'd11, 3'd0}, {6'd12, 3'd0}, {6'd13, 3'd0}:
            Alphabet = 5'd9;
        {6'd11, 3'd1}, {6'd11, 3'd2}, {6'd11, 3'd3}, {6'd11, 3'd4}, {6'd11, 3'd5},
        {6'd12, 3'd1}, {6'd12, 3'd2}, {6'd12, 3'd3}, {6'd12, 3'd4}, {6'd12, 3'd5},
        {6'd13, 3'd1}, {6'd13, 3'd2}, {6'd13, 3'd3}, {6'd13, 3'd4}, {6'd13, 3'd5}:
            Alphabet = 5'd10;

        default: Alphabet = 5'd0;
    endcase
end

endmodule
